`default_nettype none

// TODO implement signature export as required by RISCOF before finish is
// called

module control #(
    parameter integer BASE_ADDRESS
) (
    input wire clk_i,
    input wire rst_i,
    input wire stb_i,
    input wire cyc_i,
    input wire[31:0] adr_i,
    input wire[3:0] sel_i,
    input wire[31:0] dat_i,
    output reg[31:0] dat_o,
    input wire we_i,
    output reg ack_o,
    output reg err_o,
    output reg rty_o
);

always @(posedge clk_i) begin
    ack_o <= 0;
    err_o <= 0;
    rty_o <= 0;
    dat_o <= 32'hzzzz_zzzz;

    if (stb_i & cyc_i & adr_i == BASE_ADDRESS) begin
        $display("Control register accessed, finishing simulation");
        $finish;
    end
end

endmodule

`default_nettype none

module alu(
   input wire[0:31] instruction;
);



endmodule

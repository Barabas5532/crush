`default_nettype none

module alu_tb();

initial
  begin
    $display("Hello World!");
    $finish ;
  end

endmodule
